interface full_adder_if;
  logic a;
  logic b;
  logic c;
  logic sum;
  logic carry;
endinterface